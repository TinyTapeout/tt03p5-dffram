module RAM32 (CLK,
    EN0,
    VGND,
    VPWR,
    A0,
    Di0,
    Do0,
    WE0);
 input CLK;
 input EN0;
 input VGND;
 input VPWR;
 input [4:0] A0;
 input [31:0] Di0;
 output [31:0] Do0;
 input [3:0] WE0;

 wire \A0BUF[0].X ;
 wire \A0BUF[1].X ;
 wire \A0BUF[2].X ;
 wire \A0BUF[3].X ;
 wire \A0BUF[4].X ;
 wire \DEC0.EN ;
 wire \DIBUF[0].X ;
 wire \DIBUF[10].X ;
 wire \DIBUF[11].X ;
 wire \DIBUF[12].X ;
 wire \DIBUF[13].X ;
 wire \DIBUF[14].X ;
 wire \DIBUF[15].X ;
 wire \DIBUF[16].X ;
 wire \DIBUF[17].X ;
 wire \DIBUF[18].X ;
 wire \DIBUF[19].X ;
 wire \DIBUF[1].X ;
 wire \DIBUF[20].X ;
 wire \DIBUF[21].X ;
 wire \DIBUF[22].X ;
 wire \DIBUF[23].X ;
 wire \DIBUF[24].X ;
 wire \DIBUF[25].X ;
 wire \DIBUF[26].X ;
 wire \DIBUF[27].X ;
 wire \DIBUF[28].X ;
 wire \DIBUF[29].X ;
 wire \DIBUF[2].X ;
 wire \DIBUF[30].X ;
 wire \DIBUF[31].X ;
 wire \DIBUF[3].X ;
 wire \DIBUF[4].X ;
 wire \DIBUF[5].X ;
 wire \DIBUF[6].X ;
 wire \DIBUF[7].X ;
 wire \DIBUF[8].X ;
 wire \DIBUF[9].X ;
 wire \Do0MUX.A0[0] ;
 wire \Do0MUX.A0[10] ;
 wire \Do0MUX.A0[11] ;
 wire \Do0MUX.A0[12] ;
 wire \Do0MUX.A0[13] ;
 wire \Do0MUX.A0[14] ;
 wire \Do0MUX.A0[15] ;
 wire \Do0MUX.A0[16] ;
 wire \Do0MUX.A0[17] ;
 wire \Do0MUX.A0[18] ;
 wire \Do0MUX.A0[19] ;
 wire \Do0MUX.A0[1] ;
 wire \Do0MUX.A0[20] ;
 wire \Do0MUX.A0[21] ;
 wire \Do0MUX.A0[22] ;
 wire \Do0MUX.A0[23] ;
 wire \Do0MUX.A0[24] ;
 wire \Do0MUX.A0[25] ;
 wire \Do0MUX.A0[26] ;
 wire \Do0MUX.A0[27] ;
 wire \Do0MUX.A0[28] ;
 wire \Do0MUX.A0[29] ;
 wire \Do0MUX.A0[2] ;
 wire \Do0MUX.A0[30] ;
 wire \Do0MUX.A0[31] ;
 wire \Do0MUX.A0[3] ;
 wire \Do0MUX.A0[4] ;
 wire \Do0MUX.A0[5] ;
 wire \Do0MUX.A0[6] ;
 wire \Do0MUX.A0[7] ;
 wire \Do0MUX.A0[8] ;
 wire \Do0MUX.A0[9] ;
 wire \Do0MUX.A1[0] ;
 wire \Do0MUX.A1[10] ;
 wire \Do0MUX.A1[11] ;
 wire \Do0MUX.A1[12] ;
 wire \Do0MUX.A1[13] ;
 wire \Do0MUX.A1[14] ;
 wire \Do0MUX.A1[15] ;
 wire \Do0MUX.A1[16] ;
 wire \Do0MUX.A1[17] ;
 wire \Do0MUX.A1[18] ;
 wire \Do0MUX.A1[19] ;
 wire \Do0MUX.A1[1] ;
 wire \Do0MUX.A1[20] ;
 wire \Do0MUX.A1[21] ;
 wire \Do0MUX.A1[22] ;
 wire \Do0MUX.A1[23] ;
 wire \Do0MUX.A1[24] ;
 wire \Do0MUX.A1[25] ;
 wire \Do0MUX.A1[26] ;
 wire \Do0MUX.A1[27] ;
 wire \Do0MUX.A1[28] ;
 wire \Do0MUX.A1[29] ;
 wire \Do0MUX.A1[2] ;
 wire \Do0MUX.A1[30] ;
 wire \Do0MUX.A1[31] ;
 wire \Do0MUX.A1[3] ;
 wire \Do0MUX.A1[4] ;
 wire \Do0MUX.A1[5] ;
 wire \Do0MUX.A1[6] ;
 wire \Do0MUX.A1[7] ;
 wire \Do0MUX.A1[8] ;
 wire \Do0MUX.A1[9] ;
 wire \Do0MUX.SEL[0] ;
 wire \Do0MUX.SEL[1] ;
 wire \Do0MUX.SEL[2] ;
 wire \Do0MUX.SEL[3] ;
 wire \SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ;
 wire \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ;
 wire \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ;
 wire \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ;
 wire \SLICE_16[0].RAM16.CLKBUF.X ;
 wire \SLICE_16[0].RAM16.DEC0.EN ;
 wire \SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ;
 wire \SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ;
 wire \SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ;
 wire \SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ;
 wire \SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \SLICE_16[0].RAM16.EN0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].A ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].A ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].A ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].A ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE_16[0].RAM16.WEBUF[0].A ;
 wire \SLICE_16[0].RAM16.WEBUF[1].A ;
 wire \SLICE_16[0].RAM16.WEBUF[2].A ;
 wire \SLICE_16[0].RAM16.WEBUF[3].A ;
 wire \SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ;
 wire \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ;
 wire \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ;
 wire \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ;
 wire \SLICE_16[1].RAM16.CLKBUF.X ;
 wire \SLICE_16[1].RAM16.DEC0.EN ;
 wire \SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ;
 wire \SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ;
 wire \SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ;
 wire \SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ;
 wire \SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \SLICE_16[1].RAM16.EN0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].A ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].A ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].A ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].A ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;

 sky130_fd_sc_hd__clkbuf_2 \A0BUF[0].__cell__  (.A(A0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[1].__cell__  (.A(A0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[2].__cell__  (.A(A0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[3].__cell__  (.A(A0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[4].__cell__  (.A(A0[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \DEC0.AND0  (.A_N(\A0BUF[4].X ),
    .B(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \DEC0.AND1  (.A(\A0BUF[4].X ),
    .B(\DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[0].__cell__  (.A(Di0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[10].__cell__  (.A(Di0[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[11].__cell__  (.A(Di0[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[12].__cell__  (.A(Di0[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[13].__cell__  (.A(Di0[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[14].__cell__  (.A(Di0[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[15].__cell__  (.A(Di0[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[16].__cell__  (.A(Di0[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[17].__cell__  (.A(Di0[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[18].__cell__  (.A(Di0[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[19].__cell__  (.A(Di0[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[1].__cell__  (.A(Di0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[20].__cell__  (.A(Di0[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[21].__cell__  (.A(Di0[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[22].__cell__  (.A(Di0[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[23].__cell__  (.A(Di0[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[24].__cell__  (.A(Di0[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[25].__cell__  (.A(Di0[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[26].__cell__  (.A(Di0[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[27].__cell__  (.A(Di0[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[28].__cell__  (.A(Di0[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[29].__cell__  (.A(Di0[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[2].__cell__  (.A(Di0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[30].__cell__  (.A(Di0[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[31].__cell__  (.A(Di0[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[3].__cell__  (.A(Di0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[4].__cell__  (.A(Di0[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[5].__cell__  (.A(Di0[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[6].__cell__  (.A(Di0[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[7].__cell__  (.A(Di0[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[8].__cell__  (.A(Di0[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[9].__cell__  (.A(Di0[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DIBUF[9].X ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\Do0MUX.A0[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\Do0MUX.A0[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\Do0MUX.A0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\Do0MUX.A0[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\Do0MUX.A0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\Do0MUX.A0[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\Do0MUX.A0[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\Do0MUX.A0[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\Do0MUX.A1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\Do0MUX.A1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\Do0MUX.A1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\Do0MUX.A1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\Do0MUX.A1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\Do0MUX.A1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\Do0MUX.A1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\Do0MUX.A1[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[0]  (.A0(\Do0MUX.A0[0] ),
    .A1(\Do0MUX.A1[0] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[0]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[1]  (.A0(\Do0MUX.A0[1] ),
    .A1(\Do0MUX.A1[1] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[1]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[2]  (.A0(\Do0MUX.A0[2] ),
    .A1(\Do0MUX.A1[2] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[2]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[3]  (.A0(\Do0MUX.A0[3] ),
    .A1(\Do0MUX.A1[3] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[3]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[4]  (.A0(\Do0MUX.A0[4] ),
    .A1(\Do0MUX.A1[4] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[4]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[5]  (.A0(\Do0MUX.A0[5] ),
    .A1(\Do0MUX.A1[5] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[5]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[6]  (.A0(\Do0MUX.A0[6] ),
    .A1(\Do0MUX.A1[6] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[6]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[7]  (.A0(\Do0MUX.A0[7] ),
    .A1(\Do0MUX.A1[7] ),
    .S(\Do0MUX.SEL[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[7]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[10]  (.DIODE(\Do0MUX.A0[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[11]  (.DIODE(\Do0MUX.A0[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[12]  (.DIODE(\Do0MUX.A0[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[13]  (.DIODE(\Do0MUX.A0[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[14]  (.DIODE(\Do0MUX.A0[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[15]  (.DIODE(\Do0MUX.A0[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[8]  (.DIODE(\Do0MUX.A0[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[9]  (.DIODE(\Do0MUX.A0[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[10]  (.DIODE(\Do0MUX.A1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[11]  (.DIODE(\Do0MUX.A1[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[12]  (.DIODE(\Do0MUX.A1[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[13]  (.DIODE(\Do0MUX.A1[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[14]  (.DIODE(\Do0MUX.A1[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[15]  (.DIODE(\Do0MUX.A1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[8]  (.DIODE(\Do0MUX.A1[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[9]  (.DIODE(\Do0MUX.A1[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[0]  (.A0(\Do0MUX.A0[8] ),
    .A1(\Do0MUX.A1[8] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[8]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[1]  (.A0(\Do0MUX.A0[9] ),
    .A1(\Do0MUX.A1[9] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[9]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[2]  (.A0(\Do0MUX.A0[10] ),
    .A1(\Do0MUX.A1[10] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[10]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[3]  (.A0(\Do0MUX.A0[11] ),
    .A1(\Do0MUX.A1[11] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[11]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[4]  (.A0(\Do0MUX.A0[12] ),
    .A1(\Do0MUX.A1[12] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[12]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[5]  (.A0(\Do0MUX.A0[13] ),
    .A1(\Do0MUX.A1[13] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[13]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[6]  (.A0(\Do0MUX.A0[14] ),
    .A1(\Do0MUX.A1[14] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[14]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[1].MUX[7]  (.A0(\Do0MUX.A0[15] ),
    .A1(\Do0MUX.A1[15] ),
    .S(\Do0MUX.SEL[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[15]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[16]  (.DIODE(\Do0MUX.A0[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[17]  (.DIODE(\Do0MUX.A0[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[18]  (.DIODE(\Do0MUX.A0[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[19]  (.DIODE(\Do0MUX.A0[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[20]  (.DIODE(\Do0MUX.A0[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[21]  (.DIODE(\Do0MUX.A0[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[22]  (.DIODE(\Do0MUX.A0[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[23]  (.DIODE(\Do0MUX.A0[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[16]  (.DIODE(\Do0MUX.A1[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[17]  (.DIODE(\Do0MUX.A1[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[18]  (.DIODE(\Do0MUX.A1[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[19]  (.DIODE(\Do0MUX.A1[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[20]  (.DIODE(\Do0MUX.A1[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[21]  (.DIODE(\Do0MUX.A1[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[22]  (.DIODE(\Do0MUX.A1[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[23]  (.DIODE(\Do0MUX.A1[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[0]  (.A0(\Do0MUX.A0[16] ),
    .A1(\Do0MUX.A1[16] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[16]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[1]  (.A0(\Do0MUX.A0[17] ),
    .A1(\Do0MUX.A1[17] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[17]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[2]  (.A0(\Do0MUX.A0[18] ),
    .A1(\Do0MUX.A1[18] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[18]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[3]  (.A0(\Do0MUX.A0[19] ),
    .A1(\Do0MUX.A1[19] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[19]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[4]  (.A0(\Do0MUX.A0[20] ),
    .A1(\Do0MUX.A1[20] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[20]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[5]  (.A0(\Do0MUX.A0[21] ),
    .A1(\Do0MUX.A1[21] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[21]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[6]  (.A0(\Do0MUX.A0[22] ),
    .A1(\Do0MUX.A1[22] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[22]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[2].MUX[7]  (.A0(\Do0MUX.A0[23] ),
    .A1(\Do0MUX.A1[23] ),
    .S(\Do0MUX.SEL[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[23]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[24]  (.DIODE(\Do0MUX.A0[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[25]  (.DIODE(\Do0MUX.A0[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[26]  (.DIODE(\Do0MUX.A0[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[27]  (.DIODE(\Do0MUX.A0[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[28]  (.DIODE(\Do0MUX.A0[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[29]  (.DIODE(\Do0MUX.A0[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[30]  (.DIODE(\Do0MUX.A0[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[31]  (.DIODE(\Do0MUX.A0[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[24]  (.DIODE(\Do0MUX.A1[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[25]  (.DIODE(\Do0MUX.A1[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[26]  (.DIODE(\Do0MUX.A1[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[27]  (.DIODE(\Do0MUX.A1[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[28]  (.DIODE(\Do0MUX.A1[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[29]  (.DIODE(\Do0MUX.A1[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[30]  (.DIODE(\Do0MUX.A1[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[31]  (.DIODE(\Do0MUX.A1[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[0]  (.A0(\Do0MUX.A0[24] ),
    .A1(\Do0MUX.A1[24] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[24]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[1]  (.A0(\Do0MUX.A0[25] ),
    .A1(\Do0MUX.A1[25] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[25]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[2]  (.A0(\Do0MUX.A0[26] ),
    .A1(\Do0MUX.A1[26] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[26]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[3]  (.A0(\Do0MUX.A0[27] ),
    .A1(\Do0MUX.A1[27] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[27]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[4]  (.A0(\Do0MUX.A0[28] ),
    .A1(\Do0MUX.A1[28] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[28]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[5]  (.A0(\Do0MUX.A0[29] ),
    .A1(\Do0MUX.A1[29] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[29]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[6]  (.A0(\Do0MUX.A0[30] ),
    .A1(\Do0MUX.A1[30] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[30]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[3].MUX[7]  (.A0(\Do0MUX.A0[31] ),
    .A1(\Do0MUX.A1[31] ),
    .S(\Do0MUX.SEL[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Do0[31]));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[0]  (.A(\A0BUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0MUX.SEL[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[1]  (.A(\A0BUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0MUX.SEL[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[2]  (.A(\A0BUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0MUX.SEL[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[3]  (.A(\A0BUF[4].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Do0MUX.SEL[3] ));
 sky130_fd_sc_hd__clkbuf_2 \EN0BUF.__cell__  (.A(EN0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].__cell__  (.A(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(CLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\SLICE_16[0].RAM16.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \SLICE_16[0].RAM16.DEC0.AND1  (.A(\SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\SLICE_16[0].RAM16.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[1]  (.A(\SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[2]  (.A(\SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[3]  (.A(\SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[8] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[9] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[10] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[11] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[12] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[13] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[14] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[15] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[16] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[17] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[18] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[19] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[20] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[21] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[22] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[23] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[24] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[25] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[26] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[27] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[28] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[29] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[30] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\SLICE_16[0].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A0[31] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\SLICE_16[0].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\SLICE_16[0].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\SLICE_16[0].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.FBUFENBUF0[1].__cell__  (.A(\SLICE_16[0].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.FBUFENBUF0[2].__cell__  (.A(\SLICE_16[0].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.FBUFENBUF0[3].__cell__  (.A(\SLICE_16[0].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\SLICE_16[0].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\SLICE_16[0].RAM16.A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\SLICE_16[0].RAM16.A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\SLICE_16[0].RAM16.A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\SLICE_16[0].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\SLICE_16[0].RAM16.A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\SLICE_16[0].RAM16.A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\SLICE_16[0].RAM16.A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[0].RAM16.TIE0[0].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[0].RAM16.TIE0[1].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[0].RAM16.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[0].RAM16.TIE0[2].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[0].RAM16.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[0].RAM16.TIE0[3].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[0].RAM16.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.WEBUF[1].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.WEBUF[2].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[0].RAM16.WEBUF[3].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].__cell__  (.A(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(CLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\SLICE_16[1].RAM16.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \SLICE_16[1].RAM16.DEC0.AND1  (.A(\SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\SLICE_16[1].RAM16.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[1]  (.A(\SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[2]  (.A(\SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[3]  (.A(\SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[0] ),
    .D(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[7] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[8] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[9] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[10] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[11] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[12] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[13] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[14] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[1] ),
    .D(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[15] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[16] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[17] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[18] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[19] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[20] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[21] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[22] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[2] ),
    .D(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[23] ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[24] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[25] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[26] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[27] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[28] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[29] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[30] ));
 sky130_fd_sc_hd__dfxtp_1 \SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\SLICE_16[1].RAM16.Do0_REG.CLKBUF[3] ),
    .D(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Do0MUX.A1[31] ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\SLICE_16[1].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\SLICE_16[1].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\SLICE_16[1].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.FBUFENBUF0[1].__cell__  (.A(\SLICE_16[1].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.FBUFENBUF0[2].__cell__  (.A(\SLICE_16[1].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.FBUFENBUF0[3].__cell__  (.A(\SLICE_16[1].RAM16.EN0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\SLICE_16[1].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\SLICE_16[1].RAM16.A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\SLICE_16[1].RAM16.A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\SLICE_16[1].RAM16.A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\SLICE_16[1].RAM16.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\SLICE_16[1].RAM16.A0BUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\SLICE_16[1].RAM16.A0BUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\SLICE_16[1].RAM16.A0BUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[1].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[2].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[3].X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .GCLK(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[1].RAM16.TIE0[0].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[1].RAM16.TIE0[1].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[1].RAM16.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[1].RAM16.TIE0[2].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[1].RAM16.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \SLICE_16[1].RAM16.TIE0[3].__cell__  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(\SLICE_16[1].RAM16.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[0].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.WEBUF[1].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[1].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.WEBUF[2].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[2].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \SLICE_16[1].RAM16.WEBUF[3].__cell__  (.A(\SLICE_16[0].RAM16.WEBUF[3].A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[0].__cell__  (.A(WE0[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[1].__cell__  (.A(WE0[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[2].__cell__  (.A(WE0[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[3].__cell__  (.A(WE0[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SLICE_16[0].RAM16.WEBUF[3].A ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_0_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_0_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_10_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_10_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_11_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_12_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_12_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_13_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_13_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_13_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_14_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_14_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_14_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_14_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_15_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_15_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_15_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_16_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_16_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_16_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_16_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_17_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_17_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_17_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_17_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_17_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_18_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_18_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_18_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_20_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_22_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_22_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_22_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_23_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_23_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_23_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_24_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_24_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_24_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_24_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_25_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_25_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_25_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_26_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_26_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_26_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_26_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_28_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_28_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_29_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_2_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_30_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_30_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_31_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_31_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_31_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_32_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_32_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_32_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_32_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_33_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_33_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_33_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_34_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_34_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_34_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_34_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_35_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_35_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_35_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_35_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_35_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 fill_36_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_36_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_36_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_36_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_37_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_37_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_77 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_37_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_37_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_38_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 fill_38_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_3_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_4_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_4_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_4_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 fill_5_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_5_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_5_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_6_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_6_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_6_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_6_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_7_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_7_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 fill_8_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_8_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_8_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 fill_8_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 fill_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_0 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_1 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_11 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_16 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_17 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_18 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_19 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_2 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_20 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_21 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_22 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_23 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_24 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_25 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_26 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_27 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_28 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_29 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_3 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_4 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_5 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_9 (.VGND(VGND),
    .VPWR(VPWR));
endmodule
