module RAM32(
  input CLK,
  input [4:0] A0,
  input [3:0] WE0,
  input EN0,
  input [31:0] Di0,
  output [31:0] Do0
);

endmodule
