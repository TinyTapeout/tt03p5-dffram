VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 401.580 BY 111.520 ;
  PIN A0[0]
    PORT
      LAYER met3 ;
        RECT 399.580 16.360 401.580 16.960 ;
    END
  END A0[0]
  PIN A0[1]
    PORT
      LAYER met3 ;
        RECT 399.580 25.880 401.580 26.480 ;
    END
  END A0[1]
  PIN A0[2]
    PORT
      LAYER met3 ;
        RECT 399.580 35.400 401.580 36.000 ;
    END
  END A0[2]
  PIN A0[3]
    PORT
      LAYER met3 ;
        RECT 399.580 44.920 401.580 45.520 ;
    END
  END A0[3]
  PIN A0[4]
    PORT
      LAYER met3 ;
        RECT 399.580 54.440 401.580 55.040 ;
    END
  END A0[4]
  PIN CLK
    PORT
      LAYER met3 ;
        RECT 399.580 63.960 401.580 64.560 ;
    END
  END CLK
  PIN Di0[0]
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    PORT
      LAYER met2 ;
        RECT 7.910 109.520 8.190 111.520 ;
    END
  END Do0[0]
  PIN Do0[10]
    PORT
      LAYER met2 ;
        RECT 132.110 109.520 132.390 111.520 ;
    END
  END Do0[10]
  PIN Do0[11]
    PORT
      LAYER met2 ;
        RECT 144.530 109.520 144.810 111.520 ;
    END
  END Do0[11]
  PIN Do0[12]
    PORT
      LAYER met2 ;
        RECT 156.950 109.520 157.230 111.520 ;
    END
  END Do0[12]
  PIN Do0[13]
    PORT
      LAYER met2 ;
        RECT 169.370 109.520 169.650 111.520 ;
    END
  END Do0[13]
  PIN Do0[14]
    PORT
      LAYER met2 ;
        RECT 181.790 109.520 182.070 111.520 ;
    END
  END Do0[14]
  PIN Do0[15]
    PORT
      LAYER met2 ;
        RECT 194.210 109.520 194.490 111.520 ;
    END
  END Do0[15]
  PIN Do0[16]
    PORT
      LAYER met2 ;
        RECT 206.630 109.520 206.910 111.520 ;
    END
  END Do0[16]
  PIN Do0[17]
    PORT
      LAYER met2 ;
        RECT 219.050 109.520 219.330 111.520 ;
    END
  END Do0[17]
  PIN Do0[18]
    PORT
      LAYER met2 ;
        RECT 231.470 109.520 231.750 111.520 ;
    END
  END Do0[18]
  PIN Do0[19]
    PORT
      LAYER met2 ;
        RECT 243.890 109.520 244.170 111.520 ;
    END
  END Do0[19]
  PIN Do0[1]
    PORT
      LAYER met2 ;
        RECT 20.330 109.520 20.610 111.520 ;
    END
  END Do0[1]
  PIN Do0[20]
    PORT
      LAYER met2 ;
        RECT 256.310 109.520 256.590 111.520 ;
    END
  END Do0[20]
  PIN Do0[21]
    PORT
      LAYER met2 ;
        RECT 268.730 109.520 269.010 111.520 ;
    END
  END Do0[21]
  PIN Do0[22]
    PORT
      LAYER met2 ;
        RECT 281.150 109.520 281.430 111.520 ;
    END
  END Do0[22]
  PIN Do0[23]
    PORT
      LAYER met2 ;
        RECT 293.570 109.520 293.850 111.520 ;
    END
  END Do0[23]
  PIN Do0[24]
    PORT
      LAYER met2 ;
        RECT 305.990 109.520 306.270 111.520 ;
    END
  END Do0[24]
  PIN Do0[25]
    PORT
      LAYER met2 ;
        RECT 318.410 109.520 318.690 111.520 ;
    END
  END Do0[25]
  PIN Do0[26]
    PORT
      LAYER met2 ;
        RECT 330.830 109.520 331.110 111.520 ;
    END
  END Do0[26]
  PIN Do0[27]
    PORT
      LAYER met2 ;
        RECT 343.250 109.520 343.530 111.520 ;
    END
  END Do0[27]
  PIN Do0[28]
    PORT
      LAYER met2 ;
        RECT 355.670 109.520 355.950 111.520 ;
    END
  END Do0[28]
  PIN Do0[29]
    PORT
      LAYER met2 ;
        RECT 368.090 109.520 368.370 111.520 ;
    END
  END Do0[29]
  PIN Do0[2]
    PORT
      LAYER met2 ;
        RECT 32.750 109.520 33.030 111.520 ;
    END
  END Do0[2]
  PIN Do0[30]
    PORT
      LAYER met2 ;
        RECT 380.510 109.520 380.790 111.520 ;
    END
  END Do0[30]
  PIN Do0[31]
    PORT
      LAYER met2 ;
        RECT 392.930 109.520 393.210 111.520 ;
    END
  END Do0[31]
  PIN Do0[3]
    PORT
      LAYER met2 ;
        RECT 45.170 109.520 45.450 111.520 ;
    END
  END Do0[3]
  PIN Do0[4]
    PORT
      LAYER met2 ;
        RECT 57.590 109.520 57.870 111.520 ;
    END
  END Do0[4]
  PIN Do0[5]
    PORT
      LAYER met2 ;
        RECT 70.010 109.520 70.290 111.520 ;
    END
  END Do0[5]
  PIN Do0[6]
    PORT
      LAYER met2 ;
        RECT 82.430 109.520 82.710 111.520 ;
    END
  END Do0[6]
  PIN Do0[7]
    PORT
      LAYER met2 ;
        RECT 94.850 109.520 95.130 111.520 ;
    END
  END Do0[7]
  PIN Do0[8]
    PORT
      LAYER met2 ;
        RECT 107.270 109.520 107.550 111.520 ;
    END
  END Do0[8]
  PIN Do0[9]
    PORT
      LAYER met2 ;
        RECT 119.690 109.520 119.970 111.520 ;
    END
  END Do0[9]
  PIN EN0
    PORT
      LAYER met3 ;
        RECT 399.580 6.840 401.580 7.440 ;
    END
  END EN0
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 109.040 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 109.040 ;
    END
  END VPWR
  PIN WE0[0]
    PORT
      LAYER met3 ;
        RECT 399.580 73.480 401.580 74.080 ;
    END
  END WE0[0]
  PIN WE0[1]
    PORT
      LAYER met3 ;
        RECT 399.580 83.000 401.580 83.600 ;
    END
  END WE0[1]
  PIN WE0[2]
    PORT
      LAYER met3 ;
        RECT 399.580 92.520 401.580 93.120 ;
    END
  END WE0[2]
  PIN WE0[3]
    PORT
      LAYER met3 ;
        RECT 399.580 102.040 401.580 102.640 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 399.010 108.990 ;
        RECT 2.570 101.945 399.010 104.775 ;
        RECT 2.570 96.555 399.010 99.335 ;
        RECT 2.570 96.505 84.715 96.555 ;
        RECT 2.570 93.845 85.175 93.895 ;
        RECT 2.570 91.115 399.010 93.845 ;
        RECT 2.570 91.065 84.715 91.115 ;
        RECT 2.570 88.405 85.175 88.455 ;
        RECT 2.570 85.675 399.010 88.405 ;
        RECT 2.570 85.625 84.715 85.675 ;
        RECT 2.570 82.965 85.175 83.015 ;
        RECT 2.570 80.235 399.010 82.965 ;
        RECT 2.570 80.185 84.715 80.235 ;
        RECT 2.570 77.525 85.175 77.575 ;
        RECT 2.570 74.795 399.010 77.525 ;
        RECT 2.570 74.745 84.715 74.795 ;
        RECT 2.570 72.085 85.175 72.135 ;
        RECT 2.570 69.355 399.010 72.085 ;
        RECT 2.570 69.305 84.715 69.355 ;
        RECT 2.570 66.645 85.175 66.695 ;
        RECT 2.570 63.915 399.010 66.645 ;
        RECT 2.570 63.865 84.715 63.915 ;
        RECT 2.570 61.205 85.175 61.255 ;
        RECT 2.570 58.475 399.010 61.205 ;
        RECT 2.570 58.425 84.715 58.475 ;
        RECT 2.570 55.765 85.175 55.815 ;
        RECT 2.570 52.985 399.010 55.765 ;
        RECT 2.570 47.595 399.010 50.375 ;
        RECT 2.570 47.545 84.715 47.595 ;
        RECT 2.570 44.885 85.175 44.935 ;
        RECT 2.570 42.155 399.010 44.885 ;
        RECT 2.570 42.105 84.715 42.155 ;
        RECT 2.570 39.445 85.175 39.495 ;
        RECT 2.570 36.715 399.010 39.445 ;
        RECT 2.570 36.665 84.715 36.715 ;
        RECT 2.570 34.005 85.175 34.055 ;
        RECT 2.570 31.275 399.010 34.005 ;
        RECT 2.570 31.225 84.715 31.275 ;
        RECT 2.570 28.565 85.175 28.615 ;
        RECT 2.570 25.835 399.010 28.565 ;
        RECT 2.570 25.785 84.715 25.835 ;
        RECT 2.570 23.125 85.175 23.175 ;
        RECT 2.570 20.395 399.010 23.125 ;
        RECT 2.570 20.345 84.715 20.395 ;
        RECT 2.570 17.685 85.175 17.735 ;
        RECT 2.570 14.955 399.010 17.685 ;
        RECT 2.570 14.905 84.715 14.955 ;
        RECT 2.570 12.245 85.175 12.295 ;
        RECT 2.570 9.515 399.010 12.245 ;
        RECT 2.570 9.465 84.715 9.515 ;
        RECT 2.570 6.805 85.175 6.855 ;
        RECT 2.570 4.025 399.010 6.805 ;
      LAYER li1 ;
        RECT 2.760 2.635 398.820 108.885 ;
      LAYER met1 ;
        RECT 2.760 0.040 399.210 111.480 ;
      LAYER met2 ;
        RECT 3.310 109.240 7.630 111.510 ;
        RECT 8.470 109.240 20.050 111.510 ;
        RECT 20.890 109.240 32.470 111.510 ;
        RECT 33.310 109.240 44.890 111.510 ;
        RECT 45.730 109.240 57.310 111.510 ;
        RECT 58.150 109.240 69.730 111.510 ;
        RECT 70.570 109.240 82.150 111.510 ;
        RECT 82.990 109.240 94.570 111.510 ;
        RECT 95.410 109.240 106.990 111.510 ;
        RECT 107.830 109.240 119.410 111.510 ;
        RECT 120.250 109.240 131.830 111.510 ;
        RECT 132.670 109.240 144.250 111.510 ;
        RECT 145.090 109.240 156.670 111.510 ;
        RECT 157.510 109.240 169.090 111.510 ;
        RECT 169.930 109.240 181.510 111.510 ;
        RECT 182.350 109.240 193.930 111.510 ;
        RECT 194.770 109.240 206.350 111.510 ;
        RECT 207.190 109.240 218.770 111.510 ;
        RECT 219.610 109.240 231.190 111.510 ;
        RECT 232.030 109.240 243.610 111.510 ;
        RECT 244.450 109.240 256.030 111.510 ;
        RECT 256.870 109.240 268.450 111.510 ;
        RECT 269.290 109.240 280.870 111.510 ;
        RECT 281.710 109.240 293.290 111.510 ;
        RECT 294.130 109.240 305.710 111.510 ;
        RECT 306.550 109.240 318.130 111.510 ;
        RECT 318.970 109.240 330.550 111.510 ;
        RECT 331.390 109.240 342.970 111.510 ;
        RECT 343.810 109.240 355.390 111.510 ;
        RECT 356.230 109.240 367.810 111.510 ;
        RECT 368.650 109.240 380.230 111.510 ;
        RECT 381.070 109.240 392.650 111.510 ;
        RECT 393.490 109.240 399.180 111.510 ;
        RECT 3.310 2.280 399.180 109.240 ;
        RECT 3.310 0.010 7.630 2.280 ;
        RECT 8.470 0.010 20.050 2.280 ;
        RECT 20.890 0.010 32.470 2.280 ;
        RECT 33.310 0.010 44.890 2.280 ;
        RECT 45.730 0.010 57.310 2.280 ;
        RECT 58.150 0.010 69.730 2.280 ;
        RECT 70.570 0.010 82.150 2.280 ;
        RECT 82.990 0.010 94.570 2.280 ;
        RECT 95.410 0.010 106.990 2.280 ;
        RECT 107.830 0.010 119.410 2.280 ;
        RECT 120.250 0.010 131.830 2.280 ;
        RECT 132.670 0.010 144.250 2.280 ;
        RECT 145.090 0.010 156.670 2.280 ;
        RECT 157.510 0.010 169.090 2.280 ;
        RECT 169.930 0.010 181.510 2.280 ;
        RECT 182.350 0.010 193.930 2.280 ;
        RECT 194.770 0.010 206.350 2.280 ;
        RECT 207.190 0.010 218.770 2.280 ;
        RECT 219.610 0.010 231.190 2.280 ;
        RECT 232.030 0.010 243.610 2.280 ;
        RECT 244.450 0.010 256.030 2.280 ;
        RECT 256.870 0.010 268.450 2.280 ;
        RECT 269.290 0.010 280.870 2.280 ;
        RECT 281.710 0.010 293.290 2.280 ;
        RECT 294.130 0.010 305.710 2.280 ;
        RECT 306.550 0.010 318.130 2.280 ;
        RECT 318.970 0.010 330.550 2.280 ;
        RECT 331.390 0.010 342.970 2.280 ;
        RECT 343.810 0.010 355.390 2.280 ;
        RECT 356.230 0.010 367.810 2.280 ;
        RECT 368.650 0.010 380.230 2.280 ;
        RECT 381.070 0.010 392.650 2.280 ;
        RECT 393.490 0.010 399.180 2.280 ;
      LAYER met3 ;
        RECT 3.285 103.040 399.580 111.345 ;
        RECT 3.285 101.640 399.180 103.040 ;
        RECT 3.285 93.520 399.580 101.640 ;
        RECT 3.285 92.120 399.180 93.520 ;
        RECT 3.285 84.000 399.580 92.120 ;
        RECT 3.285 82.600 399.180 84.000 ;
        RECT 3.285 74.480 399.580 82.600 ;
        RECT 3.285 73.080 399.180 74.480 ;
        RECT 3.285 64.960 399.580 73.080 ;
        RECT 3.285 63.560 399.180 64.960 ;
        RECT 3.285 55.440 399.580 63.560 ;
        RECT 3.285 54.040 399.180 55.440 ;
        RECT 3.285 45.920 399.580 54.040 ;
        RECT 3.285 44.520 399.180 45.920 ;
        RECT 3.285 36.400 399.580 44.520 ;
        RECT 3.285 35.000 399.180 36.400 ;
        RECT 3.285 26.880 399.580 35.000 ;
        RECT 3.285 25.480 399.180 26.880 ;
        RECT 3.285 17.360 399.580 25.480 ;
        RECT 3.285 15.960 399.180 17.360 ;
        RECT 3.285 7.840 399.580 15.960 ;
        RECT 3.285 6.440 399.180 7.840 ;
        RECT 3.285 0.175 399.580 6.440 ;
      LAYER met4 ;
        RECT 143.815 30.095 171.480 106.585 ;
        RECT 173.880 30.095 248.280 106.585 ;
        RECT 250.680 30.095 325.080 106.585 ;
        RECT 327.480 30.095 393.465 106.585 ;
  END
END RAM32
END LIBRARY

